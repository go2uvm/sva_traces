interface future_gclk_if (input clk);
   
 logic req, ack;
   clocking cb @(posedge clk);
     output    req;
    output     ack ;
   endclocking : cb
 endinterface : future_gclk_if  

 import uvm_pkg::*;
   `include "uvm_macros.svh"
 
 import vw_go2uvm_pkg::*;

 class uvm_sva_test extends go2uvm_base_test;
   virtual future_gclk_if vif;
    task reset ();
    `uvm_info(log_id, "Start of reset", UVM_MEDIUM)
    repeat(10) @ (vif.cb);
    `uvm_info(log_id, "End of reset", UVM_MEDIUM)
  endtask : reset

  task main();
     int i;
    `uvm_info(log_id, "Start of Test", UVM_MEDIUM)
          


 // initial begin : stim
    repeat(100)@ (vif.cb);

         
    {vif.req, vif.ack} <= 2'b11;
    @ (vif.cb);
    {vif.cb.req,vif.ack}<=2'b00;
      
    repeat(10) @(vif.cb);
   
    {vif.cb.req, vif.cb.ack} <= 2'b10;
     @ (vif.cb);
    {vif.cb.req, vif.cb.ack} <= 2'b01;
    @ (vif.cb);
    {vif.cb.req, vif.cb.ack} <= 2'b00;
    repeat(10) @(vif.cb);
    $finish;
  //end : stim

    `uvm_info(log_id, "End of Test", UVM_MEDIUM)
    endtask : main

endclass : uvm_sva_test

//`timescale 1ns/100
module top;
   timeunit 1ns;
   timeprecision 1ns;

  logic clk = 0;
  initial forever #10 clk = !clk;
 
  //Instantiate the Interface 
 future_gclk_if if_0 (.*);

  future_gclk_test dut (.clk(clk),
                     .req(if_0.req),
		     .ack(if_0.ack)
                    );

 uvm_sva_test test_0;

  initial begin
    test_0 = new();
    test_0.vif = if_0;
    run_test();
   end
  endmodule 
