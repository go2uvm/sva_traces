module top2;
  timeunit 1ns;
  timeprecision 1ns;
logic clk, a, b, c, rst;
  logic [7:0] [7:0] ix;
  logic [2:0]  i=3, j;

  

default clocking @(negedge clk); endclocking
int ii = 5;
  initial begin
    $display("ii=%0d", ++ii);
  end


 k dut (.*);
  
        
endmodule : top2

