module m1;
    timeunit 1ns;
    timeprecision 1ns;
    logic  clk, req, ack, done, intrpt, reset_n;
    logic hdk_err; 
   m dut (.*);

endmodule : m1
