/*
Code for use with the book
"SystemVerilog Assertions Handbook, 2nd edition"ISBN  878-0-9705394-8-7

Code is copyright of VhdlCohen Publishing & CVC Pvt Ltd., copyright 2009 

www.systemverilog.us  ben@systemverilog.us
www.cvcblr.com, info@cvcblr.com

All code provided in this book and in the accompanied website is distributed
 with *ABSOLUTELY NO SUPPORT* and *NO WARRANTY* from the authors.  Neither
the authors nor any supporting vendors shall be liable for damage in connection
with, or arising out of, the furnishing, performance or use of the models
provided in the book and website.
*/
module bit_width(input clk,load=1'b1,logic [3:0] count = 4'h0,input [3:0] prevcount); 
  timeunit 1ns;
  timeprecision 100ps;
  //logic clk = 0;
  //logic load = 1'b1;
  //logic [3:0] count = 4'h0;
  //logic [3:0] prevcount;
  wire eq_ok1, eq_ok2, eq32;
  //initial forever #20 clk = ~clk; 
  
  property OK1; @ (posedge clk)  
     load |=>   count == $past(count) + 1'b1; endproperty : OK1

  property OK2; @ (posedge clk)  
    load |=>   count == 4'($past(count) + 1); endproperty : OK2

  property BAD; 
    @ (posedge clk)   load |=>   count == $past(count) + 1;  endproperty : BAD //  L

  OK1_1 : assert property (OK1);
  OK2_1 : assert property (OK2);
  BAD_1 : assert property (BAD);

   assign eq_ok1   = (count == (prevcount + 1'b1));
  assign eq_ok2   = (count == 4'(prevcount + 1));
  assign eq32 = (count == (prevcount + 1));
endmodule : bit_width
