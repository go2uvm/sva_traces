module top2;
  timeunit 1ns;
  timeprecision 1ns;
logic w, y, clk;
  

default clocking @(negedge clk); endclocking
int i = 0,j=0 ;
 

 k dut (.*);
  
        
endmodule : top2

