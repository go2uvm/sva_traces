module m9_6(input clk,req,ack,busy,input [2:1] id=3'b000);
   // bit clk, req, ack, busy;
   // bit[2:1] id=3'b000; 
     
    ap_ReqAckBusy: assert property(@(posedge clk)$rose(req) |=>  busy s_until_with ack ); // ch9/ m9_6
    ap_ReqAckBusy2: assert property(@(posedge clk)$rose(req) |=> busy[*0:$] ##1 ack && busy); 
  
    ap_poor_format: assert property(@(posedge clk) 
$rose(req) |=>  busy throughout  $rose(req)  ##[0:$]  $rose(ack));   
    //The way it is written, req and busy are both generated by the same device
    //  (since they are active on the same clock).  

    apReqAckBusy2: assert property(@(posedge clk)$rose(req) |=> 
        busy[*0:$] ##1 $rose(ack) );
        
   
endmodule : m9_6
